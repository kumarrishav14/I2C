module hvl_top();
    import uvm_pkg::*;
    initial begin
        run_test("i2c_base_test");
    end    
endmodule